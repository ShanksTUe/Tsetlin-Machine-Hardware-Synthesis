module ROM_XIN_6 #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 6,
    parameter ROM_DEPTH  = 49
) (
    input  wire [ADDR_WIDTH-1:0] addr,
    output reg [DATA_WIDTH-1:0] data
);

    // ROM Initialization
    always @(*) begin
        case (addr)
            6'h00: data = 32'b00000000000000000000000000000000;
            6'h01: data = 32'b00000000000000000000000000000000;
            6'h02: data = 32'b00000000000000000011110000000000;
            6'h03: data = 32'b11000000000000000000001111110000;
            6'h04: data = 32'b01111111000000000000000000011111;
            6'h05: data = 32'b00000011111111000000000000000000;
            6'h06: data = 32'b00000000000111110000000000000000;
            6'h07: data = 32'b00000000000000001111000000000000;
            6'h08: data = 32'b00000000000000000000111110000000;
            6'h09: data = 32'b11110000000000000000000001111110;
            6'h0A: data = 32'b00011111100000000000000000000001;
            6'h0B: data = 32'b11000000111110000000000000000000;
            6'h0C: data = 32'b11111111000001111000000000000111;
            6'h0D: data = 32'b00001111111111100011110000000000;
            6'h0E: data = 32'b00000000111111111111101111000000;
            6'h0F: data = 32'b11000000000001110000011111111100;
            6'h10: data = 32'b11111100000000000111111111111111;
            6'h11: data = 32'b11111111100000000000001111111111;
            6'h12: data = 32'b01111111111000000000000000001111;
            6'h13: data = 32'b00000000000000000000000000000000;
            6'h14: data = 32'b00000000000000000000000000000000;
            6'h15: data = 32'b00000000000000000000000000000000;
            6'h16: data = 32'b00000000000000000000000000000000;
            6'h17: data = 32'b00000000000000000000000000000000;
            6'h18: data = 32'b11111111111111110000000000000000;
            6'h19: data = 32'b11111111111111111111111111111111;
            6'h1A: data = 32'b11000011111111111111111111111111;
            6'h1B: data = 32'b11111100000011111111111111111111;
            6'h1C: data = 32'b11111111111000000011111111111111;
            6'h1D: data = 32'b11111111111111111000000011111111;
            6'h1E: data = 32'b11111111111111111111110000000011;
            6'h1F: data = 32'b00001111111111111111111111100000;
            6'h20: data = 32'b11110000011111111111111111111111;
            6'h21: data = 32'b11111111100000011111111111111111;
            6'h22: data = 32'b11111111111111100000111111111111;
            6'h23: data = 32'b11111111111111111110000001111111;
            6'h24: data = 32'b01111111111110000011111100000111;
            6'h25: data = 32'b11000011111111110000000011111000;
            6'h26: data = 32'b00000100001111111111000000000001;
            6'h27: data = 32'b11111000000000111111111100000000;
            6'h28: data = 32'b10000000000000000011111111111000;
            6'h29: data = 32'b11111100000000000000001111111111;
            6'h2A: data = 32'b11111111111100000000000001111111;
            6'h2B: data = 32'b11111111111111111000000000011111;
            6'h2C: data = 32'b11111111111111111111111111111111;
            6'h2D: data = 32'b11111111111111111111111111111111;
            6'h2E: data = 32'b11111111111111111111111111111111;
            6'h2F: data = 32'b11111111111111111111111111111111;
            6'h30: data = 32'b11111111111111111111111111111111;
            default: data = 32'b00000000000000000000000000000000;
        endcase
    end


endmodule