    // ROM Initialization
    always @(*) begin
        case (addr)
            6'h00: data = 32'b00000000000000000000000000000000;
            6'h01: data = 32'b00000000000000000000000000000000;
            6'h02: data = 32'b00000000000000000000000000000000;
            6'h03: data = 32'b00000000000000000000000000000000;
            6'h04: data = 32'b00000000000000000000000000000000;
            6'h05: data = 32'b00000000001111111100000000000000;
            6'h06: data = 32'b00000000000011111111111000000000;
            6'h07: data = 32'b00000000000000011000000001000000;
            6'h08: data = 32'b00000000000000000001100000000000;
            6'h09: data = 32'b00000000000000000000001100000000;
            6'h0A: data = 32'b10000000000000000000000000111000;
            6'h0B: data = 32'b00011000000000000000000000000011;
            6'h0C: data = 32'b00000001110000000000000000000000;
            6'h0D: data = 32'b00000000000011100000000000000000;
            6'h0E: data = 32'b00000000000000000111000000000000;
            6'h0F: data = 32'b00000000000000000000001110000000;
            6'h10: data = 32'b11000000000000000000000000011100;
            6'h11: data = 32'b11111000000000000001000000000001;
            6'h12: data = 32'b11111110000000000000000011111111;
            6'h13: data = 32'b00000000000000000000000000000011;
            6'h14: data = 32'b00000000000000000000000000000000;
            6'h15: data = 32'b00000000000000000000000000000000;
            6'h16: data = 32'b00000000000000000000000000000000;
            6'h17: data = 32'b00000000000000000000000000000000;
            6'h18: data = 32'b11111111111111110000000000000000;
            6'h19: data = 32'b11111111111111111111111111111111;
            6'h1A: data = 32'b11111111111111111111111111111111;
            6'h1B: data = 32'b11111111111111111111111111111111;
            6'h1C: data = 32'b11111111111111111111111111111111;
            6'h1D: data = 32'b00111111111111111111111111111111;
            6'h1E: data = 32'b00000001111111111111111111000000;
            6'h1F: data = 32'b01111111101111111111111111110000;
            6'h20: data = 32'b11100111111111111111111111111110;
            6'h21: data = 32'b11111100111111111111111111111111;
            6'h22: data = 32'b11111111110001111111111111111111;
            6'h23: data = 32'b11111111111111000111111111111111;
            6'h24: data = 32'b11111111111111111110011111111111;
            6'h25: data = 32'b11111111111111111111111000111111;
            6'h26: data = 32'b10001111111111111111111111110001;
            6'h27: data = 32'b11111100011111111111111111111111;
            6'h28: data = 32'b11111111111000111111111111111111;
            6'h29: data = 32'b11101111111111100011111111111111;
            6'h2A: data = 32'b11111111000000000000011111111111;
            6'h2B: data = 32'b11111111111111000000000111111111;
            6'h2C: data = 32'b11111111111111111111111111111111;
            6'h2D: data = 32'b11111111111111111111111111111111;
            6'h2E: data = 32'b11111111111111111111111111111111;
            6'h2F: data = 32'b11111111111111111111111111111111;
            6'h30: data = 32'b11111111111111111111111111111111;
            default: data = 32'b00000000000000000000000000000000;
        endcase
    end
