    // ROM Initialization
    always @(*) begin
        case (addr)
            6'h00000: data = 32'b00000000000000000000000000000000;
            6'h00001: data = 32'b00000000000000000000000000000000;
            6'h00002: data = 32'b00000000000000000000000000000000;
            6'h00003: data = 32'b00000000000000000000000000000000;
            6'h00004: data = 32'b00011111111000000000000000000000;
            6'h00005: data = 32'b00000011111111110000000000000000;
            6'h00006: data = 32'b00000000001110000111000000000000;
            6'h00007: data = 32'b00000000000000111000000000000000;
            6'h00008: data = 32'b00000000000000000001110000000000;
            6'h00009: data = 32'b10000000000000000000000111100000;
            6'h0000A: data = 32'b00111100000000000000000000001111;
            6'h0000B: data = 32'b00000011111100000000000000000000;
            6'h0000C: data = 32'b00000001111111111100000000000000;
            6'h0000D: data = 32'b00000000011110000011110000000000;
            6'h0000E: data = 32'b00000000000011100000000000000000;
            6'h0000F: data = 32'b00000000000000011100000000000000;
            6'h00010: data = 32'b00000000000000000001110000000000;
            6'h00011: data = 32'b00000000000000000000000110000000;
            6'h00012: data = 32'b11100000001000000000000000011100;
            6'h00013: data = 32'b00001111100000100000000000000001;
            6'h00014: data = 32'b00000000011111111110000000000000;
            6'h00015: data = 32'b00000000000000001111100000000000;
            6'h00016: data = 32'b00000000000000000000000000000000;
            6'h00017: data = 32'b00000000000000000000000000000000;
            6'h00018: data = 32'b11111111111111110000000000000000;
            6'h00019: data = 32'b11111111111111111111111111111111;
            6'h0001A: data = 32'b11111111111111111111111111111111;
            6'h0001B: data = 32'b11111111111111111111111111111111;
            6'h0001C: data = 32'b11111111111111111111111111111111;
            6'h0001D: data = 32'b11111111111111111110000000011111;
            6'h0001E: data = 32'b10001111111111111111110000000000;
            6'h0001F: data = 32'b01111111111111111111111111000111;
            6'h00020: data = 32'b11100011111111111111111111111100;
            6'h00021: data = 32'b11111110000111111111111111111111;
            6'h00022: data = 32'b11111111111100000111111111111111;
            6'h00023: data = 32'b11111111111111111100001111111111;
            6'h00024: data = 32'b00111111111111111111110000001111;
            6'h00025: data = 32'b11000011111111111111111000000000;
            6'h00026: data = 32'b11111111111111111111111110000111;
            6'h00027: data = 32'b00111111111111111111111111110001;
            6'h00028: data = 32'b11100011111111111111111111111110;
            6'h00029: data = 32'b11111110011111111111111111111111;
            6'h0002A: data = 32'b11111111111000111111111111111111;
            6'h0002B: data = 32'b11111111111111100001111111011111;
            6'h0002C: data = 32'b00011111111111111111000001111101;
            6'h0002D: data = 32'b00000111111111111111111110000000;
            6'h0002E: data = 32'b11111111111111111111111111111111;
            6'h0002F: data = 32'b11111111111111111111111111111111;
            6'h00030: data = 32'b11111111111111111111111111111111;
            default: data = 32'b00000000000000000000000000000000;
        endcase
    end
